//================================================================--
// Design Unit	: lab9 (structural)
//
// File Name	: ttl.v
//
// Purpose	: implement traffic light controller
//
// Author	: Peter Walsh, Vancouver Island University
//
// Environmant	: Icarus
//-------------------------------------------------------------------
// Revision List	
// Version	Author	Date	Changes
// 1.0		PW	Sept 10 New version
// 1.1		PW	June 20 2013 review
//================================================================--

module lab9 (


...

endmodule
